--dec

LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;

ENTITY dec IS
	PORT (
		S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		CL : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END dec;

ARCHITECTURE arq OF dec IS
BEGIN
	CL(0) <= (NOT S(0)) AND (NOT S(1));
	CL(1) <= (S(0)) AND (NOT S(1));
	CL(2) <= (NOT S(0)) AND (S(1));
END arq;